`include "ShiftByNBits.v"

module divideByTen(dividend, quotient, remainder);
  input [12:0] dividend;
  output [12:0] quotient;
  output [3:0] remainder;

  
  
  endmodule

