module Decoder3to8(
input [2:0] X,
input [12:0] W0,
input [12:0] W1,
input [12:0] W2,
input [12:0] W3,
input [12:0] W4,
input [12:0] W5,
input [12:0] W6,
input [12:0] W7,
output [12:0] VALUE
);



endmodule