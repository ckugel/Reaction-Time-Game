`include "dffCustom.v"

module Register(In, Load, Clock, CLRN, Q);
  input In;
  input Load;
  input Clock;
  input CLRN;
  output Q;
  
  
  assign D = Load ? In : Q;
  dffCustom regDFF (.D(D), .Clk(Clock), .CLRN(CLRN), .Q(Q), .QN(_ignore));
  
endmodule
