`ifndef divideByTenFSM
  `define divideByTenFSM

`include "divideByTenNextStateLogic.v"
module divideByTenFSM();
  
  
  
endmodule

`endif
