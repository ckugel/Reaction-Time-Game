module divideByTenNextStateLogic(S1, S0, C, I, N1, N0);
  input S1;
  input S0;
  input I;
  input C;
  output N1;
  output N0;




endmodule
