`include "tff.v"
`include "counterComponent.v"
`include "equals50k.v"

module downClock(Enable, ClkIn, ClkOut);
  input Enable;
  output ClkIn;
  output ClkOut;

   

  endmodule
