module regfile(DATAP, DATAQ, RP, RQ, WA, LD_DATA, WR, CLK);
	output [3:0] DATAP;
	output [3:0] DATAQ;
	input [2:0] RP;
	input [2:0] RQ;
	input [2:0] WA;
	input [3:0] LD_DATA;
	input WR;
	input CLK;
	
	


endmodule